
module clrtest;
    supply1 VCC;
    supply0 GND;

    //DM words
    tri0[7:0] dm_word0,dm_word1,dm_word2,dm_word3,dm_word4,dm_word5,dm_word6,dm_word7,dm_word8,dm_word9,dm_word10,dm_word11,dm_word12,dm_word13,dm_word14,dm_word15,dm_word16,dm_word17,dm_word18,dm_word19,dm_word20,dm_word21,dm_word22,dm_word23,dm_word24,dm_word25,dm_word26,dm_word27,dm_word28,dm_word29,dm_word30,dm_word31,dm_word32,dm_word33,dm_word34,dm_word35,dm_word36,dm_word37,dm_word38,dm_word39,dm_word40,dm_word41,dm_word42,dm_word43,dm_word44,dm_word45,dm_word46,dm_word47,dm_word48,dm_word49,dm_word50,dm_word51,dm_word52,dm_word53,dm_word54,dm_word55,dm_word56,dm_word57,dm_word58,dm_word59,dm_word60,dm_word61,dm_word62,dm_word63,dm_word64,dm_word65,dm_word66,dm_word67,dm_word68,dm_word69,dm_word70,dm_word71,dm_word72,dm_word73,dm_word74,dm_word75,dm_word76,dm_word77,dm_word78,dm_word79,dm_word80,dm_word81,dm_word82,dm_word83,dm_word84,dm_word85,dm_word86,dm_word87,dm_word88,dm_word89,dm_word90,dm_word91,dm_word92,dm_word93,dm_word94,dm_word95,dm_word96,dm_word97,dm_word98,dm_word99,dm_word100,dm_word101,dm_word102,dm_word103,dm_word104,dm_word105,dm_word106,dm_word107,dm_word108,dm_word109,dm_word110,dm_word111,dm_word112,dm_word113,dm_word114,dm_word115,dm_word116,dm_word117,dm_word118,dm_word119,dm_word120,dm_word121,dm_word122,dm_word123,dm_word124,dm_word125,dm_word126,dm_word127,dm_word128,dm_word129,dm_word130,dm_word131,dm_word132,dm_word133,dm_word134,dm_word135,dm_word136,dm_word137,dm_word138,dm_word139,dm_word140,dm_word141,dm_word142,dm_word143,dm_word144,dm_word145,dm_word146,dm_word147,dm_word148,dm_word149,dm_word150,dm_word151,dm_word152,dm_word153,dm_word154,dm_word155,dm_word156,dm_word157,dm_word158,dm_word159,dm_word160,dm_word161,dm_word162,dm_word163,dm_word164,dm_word165,dm_word166,dm_word167,dm_word168,dm_word169,dm_word170,dm_word171,dm_word172,dm_word173,dm_word174,dm_word175,dm_word176,dm_word177,dm_word178,dm_word179,dm_word180,dm_word181,dm_word182,dm_word183,dm_word184,dm_word185,dm_word186,dm_word187,dm_word188,dm_word189,dm_word190,dm_word191,dm_word192,dm_word193,dm_word194,dm_word195,dm_word196,dm_word197,dm_word198,dm_word199,dm_word200,dm_word201,dm_word202,dm_word203,dm_word204,dm_word205,dm_word206,dm_word207,dm_word208,dm_word209,dm_word210,dm_word211,dm_word212,dm_word213,dm_word214,dm_word215,dm_word216,dm_word217,dm_word218,dm_word219,dm_word220,dm_word221,dm_word222,dm_word223,dm_word224,dm_word225,dm_word226,dm_word227,dm_word228,dm_word229,dm_word230,dm_word231,dm_word232,dm_word233,dm_word234,dm_word235,dm_word236,dm_word237,dm_word238,dm_word239,dm_word240,dm_word241,dm_word242,dm_word243,dm_word244,dm_word245,dm_word246,dm_word247,dm_word248,dm_word249,dm_word250,dm_word251,dm_word252,dm_word253,dm_word254,dm_word255,dm_word256,dm_word257,dm_word258,dm_word259,dm_word260,dm_word261,dm_word262,dm_word263,dm_word264,dm_word265,dm_word266,dm_word267,dm_word268,dm_word269,dm_word270,dm_word271,dm_word272,dm_word273,dm_word274,dm_word275,dm_word276,dm_word277,dm_word278,dm_word279,dm_word280,dm_word281,dm_word282,dm_word283,dm_word284,dm_word285,dm_word286,dm_word287,dm_word288,dm_word289,dm_word290,dm_word291,dm_word292,dm_word293,dm_word294,dm_word295,dm_word296,dm_word297,dm_word298,dm_word299,dm_word300,dm_word301,dm_word302,dm_word303,dm_word304,dm_word305,dm_word306,dm_word307,dm_word308,dm_word309,dm_word310,dm_word311,dm_word312,dm_word313,dm_word314,dm_word315,dm_word316,dm_word317,dm_word318,dm_word319,dm_word320,dm_word321,dm_word322,dm_word323,dm_word324,dm_word325,dm_word326,dm_word327,dm_word328,dm_word329,dm_word330,dm_word331,dm_word332,dm_word333,dm_word334,dm_word335,dm_word336,dm_word337,dm_word338,dm_word339,dm_word340,dm_word341,dm_word342,dm_word343,dm_word344,dm_word345,dm_word346,dm_word347,dm_word348,dm_word349,dm_word350,dm_word351,dm_word352,dm_word353,dm_word354,dm_word355,dm_word356,dm_word357,dm_word358,dm_word359,dm_word360,dm_word361,dm_word362,dm_word363,dm_word364,dm_word365,dm_word366,dm_word367,dm_word368,dm_word369,dm_word370,dm_word371,dm_word372,dm_word373,dm_word374,dm_word375,dm_word376,dm_word377,dm_word378,dm_word379,dm_word380,dm_word381,dm_word382,dm_word383,dm_word384,dm_word385,dm_word386,dm_word387,dm_word388,dm_word389,dm_word390,dm_word391,dm_word392,dm_word393,dm_word394,dm_word395,dm_word396,dm_word397,dm_word398,dm_word399,dm_word400,dm_word401,dm_word402,dm_word403,dm_word404,dm_word405,dm_word406,dm_word407,dm_word408,dm_word409,dm_word410,dm_word411,dm_word412,dm_word413,dm_word414,dm_word415,dm_word416,dm_word417,dm_word418,dm_word419,dm_word420,dm_word421,dm_word422,dm_word423,dm_word424,dm_word425,dm_word426,dm_word427,dm_word428,dm_word429,dm_word430,dm_word431,dm_word432,dm_word433,dm_word434,dm_word435,dm_word436,dm_word437,dm_word438,dm_word439,dm_word440,dm_word441,dm_word442,dm_word443,dm_word444,dm_word445,dm_word446,dm_word447,dm_word448,dm_word449,dm_word450,dm_word451,dm_word452,dm_word453,dm_word454,dm_word455,dm_word456,dm_word457,dm_word458,dm_word459,dm_word460,dm_word461,dm_word462,dm_word463,dm_word464,dm_word465,dm_word466,dm_word467,dm_word468,dm_word469,dm_word470,dm_word471,dm_word472,dm_word473,dm_word474,dm_word475,dm_word476,dm_word477,dm_word478,dm_word479,dm_word480,dm_word481,dm_word482,dm_word483,dm_word484,dm_word485,dm_word486,dm_word487,dm_word488,dm_word489,dm_word490,dm_word491,dm_word492,dm_word493,dm_word494,dm_word495,dm_word496,dm_word497,dm_word498,dm_word499,dm_word500,dm_word501,dm_word502,dm_word503,dm_word504,dm_word505,dm_word506,dm_word507,dm_word508,dm_word509,dm_word510,dm_word511,dm_word512,dm_word513,dm_word514,dm_word515,dm_word516,dm_word517,dm_word518,dm_word519,dm_word520,dm_word521,dm_word522,dm_word523,dm_word524,dm_word525,dm_word526,dm_word527,dm_word528,dm_word529,dm_word530,dm_word531,dm_word532,dm_word533,dm_word534,dm_word535,dm_word536,dm_word537,dm_word538,dm_word539,dm_word540,dm_word541,dm_word542,dm_word543,dm_word544,dm_word545,dm_word546,dm_word547,dm_word548,dm_word549,dm_word550,dm_word551,dm_word552,dm_word553,dm_word554,dm_word555,dm_word556,dm_word557,dm_word558,dm_word559,dm_word560,dm_word561,dm_word562,dm_word563,dm_word564,dm_word565,dm_word566,dm_word567,dm_word568,dm_word569,dm_word570,dm_word571,dm_word572,dm_word573,dm_word574,dm_word575,dm_word576,dm_word577,dm_word578,dm_word579,dm_word580,dm_word581,dm_word582,dm_word583,dm_word584,dm_word585,dm_word586,dm_word587,dm_word588,dm_word589,dm_word590,dm_word591,dm_word592,dm_word593,dm_word594,dm_word595,dm_word596,dm_word597,dm_word598,dm_word599,dm_word600,dm_word601,dm_word602,dm_word603,dm_word604,dm_word605,dm_word606,dm_word607,dm_word608,dm_word609,dm_word610,dm_word611,dm_word612,dm_word613,dm_word614,dm_word615,dm_word616,dm_word617,dm_word618,dm_word619,dm_word620,dm_word621,dm_word622,dm_word623,dm_word624,dm_word625,dm_word626,dm_word627,dm_word628,dm_word629,dm_word630,dm_word631,dm_word632,dm_word633,dm_word634,dm_word635,dm_word636,dm_word637,dm_word638,dm_word639,dm_word640,dm_word641,dm_word642,dm_word643,dm_word644,dm_word645,dm_word646,dm_word647,dm_word648,dm_word649,dm_word650,dm_word651,dm_word652,dm_word653,dm_word654,dm_word655,dm_word656,dm_word657,dm_word658,dm_word659,dm_word660,dm_word661,dm_word662,dm_word663,dm_word664,dm_word665,dm_word666,dm_word667,dm_word668,dm_word669,dm_word670,dm_word671,dm_word672,dm_word673,dm_word674,dm_word675,dm_word676,dm_word677,dm_word678,dm_word679,dm_word680,dm_word681,dm_word682,dm_word683,dm_word684,dm_word685,dm_word686,dm_word687,dm_word688,dm_word689,dm_word690,dm_word691,dm_word692,dm_word693,dm_word694,dm_word695,dm_word696,dm_word697,dm_word698,dm_word699,dm_word700,dm_word701,dm_word702,dm_word703,dm_word704,dm_word705,dm_word706,dm_word707,dm_word708,dm_word709,dm_word710,dm_word711,dm_word712,dm_word713,dm_word714,dm_word715,dm_word716,dm_word717,dm_word718,dm_word719,dm_word720,dm_word721,dm_word722,dm_word723,dm_word724,dm_word725,dm_word726,dm_word727,dm_word728,dm_word729,dm_word730,dm_word731,dm_word732,dm_word733,dm_word734,dm_word735,dm_word736,dm_word737,dm_word738,dm_word739,dm_word740,dm_word741,dm_word742,dm_word743,dm_word744,dm_word745,dm_word746,dm_word747,dm_word748,dm_word749,dm_word750,dm_word751,dm_word752,dm_word753,dm_word754,dm_word755,dm_word756,dm_word757,dm_word758,dm_word759,dm_word760,dm_word761,dm_word762,dm_word763,dm_word764,dm_word765,dm_word766,dm_word767,dm_word768,dm_word769,dm_word770,dm_word771,dm_word772,dm_word773,dm_word774,dm_word775,dm_word776,dm_word777,dm_word778,dm_word779,dm_word780,dm_word781,dm_word782,dm_word783,dm_word784,dm_word785,dm_word786,dm_word787,dm_word788,dm_word789,dm_word790,dm_word791,dm_word792,dm_word793,dm_word794,dm_word795,dm_word796,dm_word797,dm_word798,dm_word799,dm_word800,dm_word801,dm_word802,dm_word803,dm_word804,dm_word805,dm_word806,dm_word807,dm_word808,dm_word809,dm_word810,dm_word811,dm_word812,dm_word813,dm_word814,dm_word815,dm_word816,dm_word817,dm_word818,dm_word819,dm_word820,dm_word821,dm_word822,dm_word823,dm_word824,dm_word825,dm_word826,dm_word827,dm_word828,dm_word829,dm_word830,dm_word831,dm_word832,dm_word833,dm_word834,dm_word835,dm_word836,dm_word837,dm_word838,dm_word839,dm_word840,dm_word841,dm_word842,dm_word843,dm_word844,dm_word845,dm_word846,dm_word847,dm_word848,dm_word849,dm_word850,dm_word851,dm_word852,dm_word853,dm_word854,dm_word855,dm_word856,dm_word857,dm_word858,dm_word859,dm_word860,dm_word861,dm_word862,dm_word863,dm_word864,dm_word865,dm_word866,dm_word867,dm_word868,dm_word869,dm_word870,dm_word871,dm_word872,dm_word873,dm_word874,dm_word875,dm_word876,dm_word877,dm_word878,dm_word879,dm_word880,dm_word881,dm_word882,dm_word883,dm_word884,dm_word885,dm_word886,dm_word887,dm_word888,dm_word889,dm_word890,dm_word891,dm_word892,dm_word893,dm_word894,dm_word895,dm_word896,dm_word897,dm_word898,dm_word899,dm_word900,dm_word901,dm_word902,dm_word903,dm_word904,dm_word905,dm_word906,dm_word907,dm_word908,dm_word909,dm_word910,dm_word911,dm_word912,dm_word913,dm_word914,dm_word915,dm_word916,dm_word917,dm_word918,dm_word919,dm_word920,dm_word921,dm_word922,dm_word923,dm_word924,dm_word925,dm_word926,dm_word927,dm_word928,dm_word929,dm_word930,dm_word931,dm_word932,dm_word933,dm_word934,dm_word935,dm_word936,dm_word937,dm_word938,dm_word939,dm_word940,dm_word941,dm_word942,dm_word943,dm_word944,dm_word945,dm_word946,dm_word947,dm_word948,dm_word949,dm_word950,dm_word951,dm_word952,dm_word953,dm_word954,dm_word955,dm_word956,dm_word957,dm_word958,dm_word959,dm_word960,dm_word961,dm_word962,dm_word963,dm_word964,dm_word965,dm_word966,dm_word967,dm_word968,dm_word969,dm_word970,dm_word971,dm_word972,dm_word973,dm_word974,dm_word975,dm_word976,dm_word977,dm_word978,dm_word979,dm_word980,dm_word981,dm_word982,dm_word983,dm_word984,dm_word985,dm_word986,dm_word987,dm_word988,dm_word989,dm_word990,dm_word991,dm_word992,dm_word993,dm_word994,dm_word995,dm_word996,dm_word997,dm_word998,dm_word999,dm_word1000,dm_word1001,dm_word1002,dm_word1003,dm_word1004,dm_word1005,dm_word1006,dm_word1007,dm_word1008,dm_word1009,dm_word1010,dm_word1011,dm_word1012,dm_word1013,dm_word1014,dm_word1015,dm_word1016,dm_word1017,dm_word1018,dm_word1019,dm_word1020,dm_word1021,dm_word1022,dm_word1023;
    //These are 'output' lines
    //PM words
    reg[15:0] pm_word0,pm_word1,pm_word2,pm_word3,pm_word4,pm_word5,pm_word6,pm_word7,pm_word8,pm_word9,pm_word10,pm_word11,pm_word12,pm_word13,pm_word14,pm_word15,pm_word16,pm_word17,pm_word18,pm_word19,pm_word20,pm_word21,pm_word22,pm_word23,pm_word24,pm_word25,pm_word26,pm_word27,pm_word28,pm_word29,pm_word30,pm_word31,pm_word32,pm_word33,pm_word34,pm_word35,pm_word36,pm_word37,pm_word38,pm_word39,pm_word40,pm_word41,pm_word42,pm_word43,pm_word44,pm_word45,pm_word46,pm_word47,pm_word48,pm_word49,pm_word50,pm_word51,pm_word52,pm_word53,pm_word54,pm_word55,pm_word56,pm_word57,pm_word58,pm_word59,pm_word60,pm_word61,pm_word62,pm_word63,pm_word64,pm_word65,pm_word66,pm_word67,pm_word68,pm_word69,pm_word70,pm_word71,pm_word72,pm_word73,pm_word74,pm_word75,pm_word76,pm_word77,pm_word78,pm_word79,pm_word80,pm_word81,pm_word82,pm_word83,pm_word84,pm_word85,pm_word86,pm_word87,pm_word88,pm_word89,pm_word90,pm_word91,pm_word92,pm_word93,pm_word94,pm_word95,pm_word96,pm_word97,pm_word98,pm_word99,pm_word100,pm_word101,pm_word102,pm_word103,pm_word104,pm_word105,pm_word106,pm_word107,pm_word108,pm_word109,pm_word110,pm_word111,pm_word112,pm_word113,pm_word114,pm_word115,pm_word116,pm_word117,pm_word118,pm_word119,pm_word120,pm_word121,pm_word122,pm_word123,pm_word124,pm_word125,pm_word126,pm_word127,pm_word128,pm_word129,pm_word130,pm_word131,pm_word132,pm_word133,pm_word134,pm_word135,pm_word136,pm_word137,pm_word138,pm_word139,pm_word140,pm_word141,pm_word142,pm_word143,pm_word144,pm_word145,pm_word146,pm_word147,pm_word148,pm_word149,pm_word150,pm_word151,pm_word152,pm_word153,pm_word154,pm_word155,pm_word156,pm_word157,pm_word158,pm_word159,pm_word160,pm_word161,pm_word162,pm_word163,pm_word164,pm_word165,pm_word166,pm_word167,pm_word168,pm_word169,pm_word170,pm_word171,pm_word172,pm_word173,pm_word174,pm_word175,pm_word176,pm_word177,pm_word178,pm_word179,pm_word180,pm_word181,pm_word182,pm_word183,pm_word184,pm_word185,pm_word186,pm_word187,pm_word188,pm_word189,pm_word190,pm_word191,pm_word192,pm_word193,pm_word194,pm_word195,pm_word196,pm_word197,pm_word198,pm_word199,pm_word200,pm_word201,pm_word202,pm_word203,pm_word204,pm_word205,pm_word206,pm_word207,pm_word208,pm_word209,pm_word210,pm_word211,pm_word212,pm_word213,pm_word214,pm_word215,pm_word216,pm_word217,pm_word218,pm_word219,pm_word220,pm_word221,pm_word222,pm_word223,pm_word224,pm_word225,pm_word226,pm_word227,pm_word228,pm_word229,pm_word230,pm_word231,pm_word232,pm_word233,pm_word234,pm_word235,pm_word236,pm_word237,pm_word238,pm_word239,pm_word240,pm_word241,pm_word242,pm_word243,pm_word244,pm_word245,pm_word246,pm_word247,pm_word248,pm_word249,pm_word250,pm_word251,pm_word252,pm_word253,pm_word254,pm_word255;
    
    reg start;                      //Active high
    tri0 clk;clock c1(clk);
    tri0[255:0] sel;                //PM sel
    tri0[1023:0] dsel;              //DM sel

    tri0[6:0] rr,r;                 //ASM enables
    tri0[4:0] rv;
    tri0[3:0] pm;
    tri0[1:0] ra,rp;
    tri0 nop,beginx;

    tri0 rd,wr;                     //Control lines-DM
    tri1 rd_latch;
    tri1 set;
    tri1 clr;

    tri0[31:26] point_add;          //Ptr- DM

    tri0 alu_write;  
    tri1[2:0] fs_cal,fs_shft;               
    tri0[7:0] alu_out,alu_flag;
    tri0 shft_wr;
    
    tri0[15:0] instruction,addbus;  //Buses
    tri0[7:0] databus;
    
    tri1[2:0] ld_val_reg;           //Control lines-PM
   
    tri0[1:0] mode;                 //PC
    
    address bu(addbus,dsel);
    datamem DM(databus,alu_out,alu_flag,dsel,point_add,clk,VCC,clr,rd,rd_latch,wr,alu_write,addbus,{dm_word1023,dm_word1022,dm_word1021,dm_word1020,dm_word1019,dm_word1018,dm_word1017,dm_word1016,dm_word1015,dm_word1014,dm_word1013,dm_word1012,dm_word1011,dm_word1010,dm_word1009,dm_word1008,dm_word1007,dm_word1006,dm_word1005,dm_word1004,dm_word1003,dm_word1002,dm_word1001,dm_word1000,dm_word999,dm_word998,dm_word997,dm_word996,dm_word995,dm_word994,dm_word993,dm_word992,dm_word991,dm_word990,dm_word989,dm_word988,dm_word987,dm_word986,dm_word985,dm_word984,dm_word983,dm_word982,dm_word981,dm_word980,dm_word979,dm_word978,dm_word977,dm_word976,dm_word975,dm_word974,dm_word973,dm_word972,dm_word971,dm_word970,dm_word969,dm_word968,dm_word967,dm_word966,dm_word965,dm_word964,dm_word963,dm_word962,dm_word961,dm_word960,dm_word959,dm_word958,dm_word957,dm_word956,dm_word955,dm_word954,dm_word953,dm_word952,dm_word951,dm_word950,dm_word949,dm_word948,dm_word947,dm_word946,dm_word945,dm_word944,dm_word943,dm_word942,dm_word941,dm_word940,dm_word939,dm_word938,dm_word937,dm_word936,dm_word935,dm_word934,dm_word933,dm_word932,dm_word931,dm_word930,dm_word929,dm_word928,dm_word927,dm_word926,dm_word925,dm_word924,dm_word923,dm_word922,dm_word921,dm_word920,dm_word919,dm_word918,dm_word917,dm_word916,dm_word915,dm_word914,dm_word913,dm_word912,dm_word911,dm_word910,dm_word909,dm_word908,dm_word907,dm_word906,dm_word905,dm_word904,dm_word903,dm_word902,dm_word901,dm_word900,dm_word899,dm_word898,dm_word897,dm_word896,dm_word895,dm_word894,dm_word893,dm_word892,dm_word891,dm_word890,dm_word889,dm_word888,dm_word887,dm_word886,dm_word885,dm_word884,dm_word883,dm_word882,dm_word881,dm_word880,dm_word879,dm_word878,dm_word877,dm_word876,dm_word875,dm_word874,dm_word873,dm_word872,dm_word871,dm_word870,dm_word869,dm_word868,dm_word867,dm_word866,dm_word865,dm_word864,dm_word863,dm_word862,dm_word861,dm_word860,dm_word859,dm_word858,dm_word857,dm_word856,dm_word855,dm_word854,dm_word853,dm_word852,dm_word851,dm_word850,dm_word849,dm_word848,dm_word847,dm_word846,dm_word845,dm_word844,dm_word843,dm_word842,dm_word841,dm_word840,dm_word839,dm_word838,dm_word837,dm_word836,dm_word835,dm_word834,dm_word833,dm_word832,dm_word831,dm_word830,dm_word829,dm_word828,dm_word827,dm_word826,dm_word825,dm_word824,dm_word823,dm_word822,dm_word821,dm_word820,dm_word819,dm_word818,dm_word817,dm_word816,dm_word815,dm_word814,dm_word813,dm_word812,dm_word811,dm_word810,dm_word809,dm_word808,dm_word807,dm_word806,dm_word805,dm_word804,dm_word803,dm_word802,dm_word801,dm_word800,dm_word799,dm_word798,dm_word797,dm_word796,dm_word795,dm_word794,dm_word793,dm_word792,dm_word791,dm_word790,dm_word789,dm_word788,dm_word787,dm_word786,dm_word785,dm_word784,dm_word783,dm_word782,dm_word781,dm_word780,dm_word779,dm_word778,dm_word777,dm_word776,dm_word775,dm_word774,dm_word773,dm_word772,dm_word771,dm_word770,dm_word769,dm_word768,dm_word767,dm_word766,dm_word765,dm_word764,dm_word763,dm_word762,dm_word761,dm_word760,dm_word759,dm_word758,dm_word757,dm_word756,dm_word755,dm_word754,dm_word753,dm_word752,dm_word751,dm_word750,dm_word749,dm_word748,dm_word747,dm_word746,dm_word745,dm_word744,dm_word743,dm_word742,dm_word741,dm_word740,dm_word739,dm_word738,dm_word737,dm_word736,dm_word735,dm_word734,dm_word733,dm_word732,dm_word731,dm_word730,dm_word729,dm_word728,dm_word727,dm_word726,dm_word725,dm_word724,dm_word723,dm_word722,dm_word721,dm_word720,dm_word719,dm_word718,dm_word717,dm_word716,dm_word715,dm_word714,dm_word713,dm_word712,dm_word711,dm_word710,dm_word709,dm_word708,dm_word707,dm_word706,dm_word705,dm_word704,dm_word703,dm_word702,dm_word701,dm_word700,dm_word699,dm_word698,dm_word697,dm_word696,dm_word695,dm_word694,dm_word693,dm_word692,dm_word691,dm_word690,dm_word689,dm_word688,dm_word687,dm_word686,dm_word685,dm_word684,dm_word683,dm_word682,dm_word681,dm_word680,dm_word679,dm_word678,dm_word677,dm_word676,dm_word675,dm_word674,dm_word673,dm_word672,dm_word671,dm_word670,dm_word669,dm_word668,dm_word667,dm_word666,dm_word665,dm_word664,dm_word663,dm_word662,dm_word661,dm_word660,dm_word659,dm_word658,dm_word657,dm_word656,dm_word655,dm_word654,dm_word653,dm_word652,dm_word651,dm_word650,dm_word649,dm_word648,dm_word647,dm_word646,dm_word645,dm_word644,dm_word643,dm_word642,dm_word641,dm_word640,dm_word639,dm_word638,dm_word637,dm_word636,dm_word635,dm_word634,dm_word633,dm_word632,dm_word631,dm_word630,dm_word629,dm_word628,dm_word627,dm_word626,dm_word625,dm_word624,dm_word623,dm_word622,dm_word621,dm_word620,dm_word619,dm_word618,dm_word617,dm_word616,dm_word615,dm_word614,dm_word613,dm_word612,dm_word611,dm_word610,dm_word609,dm_word608,dm_word607,dm_word606,dm_word605,dm_word604,dm_word603,dm_word602,dm_word601,dm_word600,dm_word599,dm_word598,dm_word597,dm_word596,dm_word595,dm_word594,dm_word593,dm_word592,dm_word591,dm_word590,dm_word589,dm_word588,dm_word587,dm_word586,dm_word585,dm_word584,dm_word583,dm_word582,dm_word581,dm_word580,dm_word579,dm_word578,dm_word577,dm_word576,dm_word575,dm_word574,dm_word573,dm_word572,dm_word571,dm_word570,dm_word569,dm_word568,dm_word567,dm_word566,dm_word565,dm_word564,dm_word563,dm_word562,dm_word561,dm_word560,dm_word559,dm_word558,dm_word557,dm_word556,dm_word555,dm_word554,dm_word553,dm_word552,dm_word551,dm_word550,dm_word549,dm_word548,dm_word547,dm_word546,dm_word545,dm_word544,dm_word543,dm_word542,dm_word541,dm_word540,dm_word539,dm_word538,dm_word537,dm_word536,dm_word535,dm_word534,dm_word533,dm_word532,dm_word531,dm_word530,dm_word529,dm_word528,dm_word527,dm_word526,dm_word525,dm_word524,dm_word523,dm_word522,dm_word521,dm_word520,dm_word519,dm_word518,dm_word517,dm_word516,dm_word515,dm_word514,dm_word513,dm_word512,dm_word511,dm_word510,dm_word509,dm_word508,dm_word507,dm_word506,dm_word505,dm_word504,dm_word503,dm_word502,dm_word501,dm_word500,dm_word499,dm_word498,dm_word497,dm_word496,dm_word495,dm_word494,dm_word493,dm_word492,dm_word491,dm_word490,dm_word489,dm_word488,dm_word487,dm_word486,dm_word485,dm_word484,dm_word483,dm_word482,dm_word481,dm_word480,dm_word479,dm_word478,dm_word477,dm_word476,dm_word475,dm_word474,dm_word473,dm_word472,dm_word471,dm_word470,dm_word469,dm_word468,dm_word467,dm_word466,dm_word465,dm_word464,dm_word463,dm_word462,dm_word461,dm_word460,dm_word459,dm_word458,dm_word457,dm_word456,dm_word455,dm_word454,dm_word453,dm_word452,dm_word451,dm_word450,dm_word449,dm_word448,dm_word447,dm_word446,dm_word445,dm_word444,dm_word443,dm_word442,dm_word441,dm_word440,dm_word439,dm_word438,dm_word437,dm_word436,dm_word435,dm_word434,dm_word433,dm_word432,dm_word431,dm_word430,dm_word429,dm_word428,dm_word427,dm_word426,dm_word425,dm_word424,dm_word423,dm_word422,dm_word421,dm_word420,dm_word419,dm_word418,dm_word417,dm_word416,dm_word415,dm_word414,dm_word413,dm_word412,dm_word411,dm_word410,dm_word409,dm_word408,dm_word407,dm_word406,dm_word405,dm_word404,dm_word403,dm_word402,dm_word401,dm_word400,dm_word399,dm_word398,dm_word397,dm_word396,dm_word395,dm_word394,dm_word393,dm_word392,dm_word391,dm_word390,dm_word389,dm_word388,dm_word387,dm_word386,dm_word385,dm_word384,dm_word383,dm_word382,dm_word381,dm_word380,dm_word379,dm_word378,dm_word377,dm_word376,dm_word375,dm_word374,dm_word373,dm_word372,dm_word371,dm_word370,dm_word369,dm_word368,dm_word367,dm_word366,dm_word365,dm_word364,dm_word363,dm_word362,dm_word361,dm_word360,dm_word359,dm_word358,dm_word357,dm_word356,dm_word355,dm_word354,dm_word353,dm_word352,dm_word351,dm_word350,dm_word349,dm_word348,dm_word347,dm_word346,dm_word345,dm_word344,dm_word343,dm_word342,dm_word341,dm_word340,dm_word339,dm_word338,dm_word337,dm_word336,dm_word335,dm_word334,dm_word333,dm_word332,dm_word331,dm_word330,dm_word329,dm_word328,dm_word327,dm_word326,dm_word325,dm_word324,dm_word323,dm_word322,dm_word321,dm_word320,dm_word319,dm_word318,dm_word317,dm_word316,dm_word315,dm_word314,dm_word313,dm_word312,dm_word311,dm_word310,dm_word309,dm_word308,dm_word307,dm_word306,dm_word305,dm_word304,dm_word303,dm_word302,dm_word301,dm_word300,dm_word299,dm_word298,dm_word297,dm_word296,dm_word295,dm_word294,dm_word293,dm_word292,dm_word291,dm_word290,dm_word289,dm_word288,dm_word287,dm_word286,dm_word285,dm_word284,dm_word283,dm_word282,dm_word281,dm_word280,dm_word279,dm_word278,dm_word277,dm_word276,dm_word275,dm_word274,dm_word273,dm_word272,dm_word271,dm_word270,dm_word269,dm_word268,dm_word267,dm_word266,dm_word265,dm_word264,dm_word263,dm_word262,dm_word261,dm_word260,dm_word259,dm_word258,dm_word257,dm_word256,dm_word255,dm_word254,dm_word253,dm_word252,dm_word251,dm_word250,dm_word249,dm_word248,dm_word247,dm_word246,dm_word245,dm_word244,dm_word243,dm_word242,dm_word241,dm_word240,dm_word239,dm_word238,dm_word237,dm_word236,dm_word235,dm_word234,dm_word233,dm_word232,dm_word231,dm_word230,dm_word229,dm_word228,dm_word227,dm_word226,dm_word225,dm_word224,dm_word223,dm_word222,dm_word221,dm_word220,dm_word219,dm_word218,dm_word217,dm_word216,dm_word215,dm_word214,dm_word213,dm_word212,dm_word211,dm_word210,dm_word209,dm_word208,dm_word207,dm_word206,dm_word205,dm_word204,dm_word203,dm_word202,dm_word201,dm_word200,dm_word199,dm_word198,dm_word197,dm_word196,dm_word195,dm_word194,dm_word193,dm_word192,dm_word191,dm_word190,dm_word189,dm_word188,dm_word187,dm_word186,dm_word185,dm_word184,dm_word183,dm_word182,dm_word181,dm_word180,dm_word179,dm_word178,dm_word177,dm_word176,dm_word175,dm_word174,dm_word173,dm_word172,dm_word171,dm_word170,dm_word169,dm_word168,dm_word167,dm_word166,dm_word165,dm_word164,dm_word163,dm_word162,dm_word161,dm_word160,dm_word159,dm_word158,dm_word157,dm_word156,dm_word155,dm_word154,dm_word153,dm_word152,dm_word151,dm_word150,dm_word149,dm_word148,dm_word147,dm_word146,dm_word145,dm_word144,dm_word143,dm_word142,dm_word141,dm_word140,dm_word139,dm_word138,dm_word137,dm_word136,dm_word135,dm_word134,dm_word133,dm_word132,dm_word131,dm_word130,dm_word129,dm_word128,dm_word127,dm_word126,dm_word125,dm_word124,dm_word123,dm_word122,dm_word121,dm_word120,dm_word119,dm_word118,dm_word117,dm_word116,dm_word115,dm_word114,dm_word113,dm_word112,dm_word111,dm_word110,dm_word109,dm_word108,dm_word107,dm_word106,dm_word105,dm_word104,dm_word103,dm_word102,dm_word101,dm_word100,dm_word99,dm_word98,dm_word97,dm_word96,dm_word95,dm_word94,dm_word93,dm_word92,dm_word91,dm_word90,dm_word89,dm_word88,dm_word87,dm_word86,dm_word85,dm_word84,dm_word83,dm_word82,dm_word81,dm_word80,dm_word79,dm_word78,dm_word77,dm_word76,dm_word75,dm_word74,dm_word73,dm_word72,dm_word71,dm_word70,dm_word69,dm_word68,dm_word67,dm_word66,dm_word65,dm_word64,dm_word63,dm_word62,dm_word61,dm_word60,dm_word59,dm_word58,dm_word57,dm_word56,dm_word55,dm_word54,dm_word53,dm_word52,dm_word51,dm_word50,dm_word49,dm_word48,dm_word47,dm_word46,dm_word45,dm_word44,dm_word43,dm_word42,dm_word41,dm_word40,dm_word39,dm_word38,dm_word37,dm_word36,dm_word35,dm_word34,dm_word33,dm_word32,dm_word31,dm_word30,dm_word29,dm_word28,dm_word27,dm_word26,dm_word25,dm_word24,dm_word23,dm_word22,dm_word21,dm_word20,dm_word19,dm_word18,dm_word17,dm_word16,dm_word15,dm_word14,dm_word13,dm_word12,dm_word11,dm_word10,dm_word9,dm_word8,dm_word7,dm_word6,dm_word5,dm_word4,dm_word3,dm_word2,dm_word1,dm_word0});
    prgrm_mem PM({pm_word255,pm_word254,pm_word253,pm_word252,pm_word251,pm_word250,pm_word249,pm_word248,pm_word247,pm_word246,pm_word245,pm_word244,pm_word243,pm_word242,pm_word241,pm_word240,pm_word239,pm_word238,pm_word237,pm_word236,pm_word235,pm_word234,pm_word233,pm_word232,pm_word231,pm_word230,pm_word229,pm_word228,pm_word227,pm_word226,pm_word225,pm_word224,pm_word223,pm_word222,pm_word221,pm_word220,pm_word219,pm_word218,pm_word217,pm_word216,pm_word215,pm_word214,pm_word213,pm_word212,pm_word211,pm_word210,pm_word209,pm_word208,pm_word207,pm_word206,pm_word205,pm_word204,pm_word203,pm_word202,pm_word201,pm_word200,pm_word199,pm_word198,pm_word197,pm_word196,pm_word195,pm_word194,pm_word193,pm_word192,pm_word191,pm_word190,pm_word189,pm_word188,pm_word187,pm_word186,pm_word185,pm_word184,pm_word183,pm_word182,pm_word181,pm_word180,pm_word179,pm_word178,pm_word177,pm_word176,pm_word175,pm_word174,pm_word173,pm_word172,pm_word171,pm_word170,pm_word169,pm_word168,pm_word167,pm_word166,pm_word165,pm_word164,pm_word163,pm_word162,pm_word161,pm_word160,pm_word159,pm_word158,pm_word157,pm_word156,pm_word155,pm_word154,pm_word153,pm_word152,pm_word151,pm_word150,pm_word149,pm_word148,pm_word147,pm_word146,pm_word145,pm_word144,pm_word143,pm_word142,pm_word141,pm_word140,pm_word139,pm_word138,pm_word137,pm_word136,pm_word135,pm_word134,pm_word133,pm_word132,pm_word131,pm_word130,pm_word129,pm_word128,pm_word127,pm_word126,pm_word125,pm_word124,pm_word123,pm_word122,pm_word121,pm_word120,pm_word119,pm_word118,pm_word117,pm_word116,pm_word115,pm_word114,pm_word113,pm_word112,pm_word111,pm_word110,pm_word109,pm_word108,pm_word107,pm_word106,pm_word105,pm_word104,pm_word103,pm_word102,pm_word101,pm_word100,pm_word99,pm_word98,pm_word97,pm_word96,pm_word95,pm_word94,pm_word93,pm_word92,pm_word91,pm_word90,pm_word89,pm_word88,pm_word87,pm_word86,pm_word85,pm_word84,pm_word83,pm_word82,pm_word81,pm_word80,pm_word79,pm_word78,pm_word77,pm_word76,pm_word75,pm_word74,pm_word73,pm_word72,pm_word71,pm_word70,pm_word69,pm_word68,pm_word67,pm_word66,pm_word65,pm_word64,pm_word63,pm_word62,pm_word61,pm_word60,pm_word59,pm_word58,pm_word57,pm_word56,pm_word55,pm_word54,pm_word53,pm_word52,pm_word51,pm_word50,pm_word49,pm_word48,pm_word47,pm_word46,pm_word45,pm_word44,pm_word43,pm_word42,pm_word41,pm_word40,pm_word39,pm_word38,pm_word37,pm_word36,pm_word35,pm_word34,pm_word33,pm_word32,pm_word31,pm_word30,pm_word29,pm_word28,pm_word27,pm_word26,pm_word25,pm_word24,pm_word23,pm_word22,pm_word21,pm_word20,pm_word19,pm_word18,pm_word17,pm_word16,pm_word15,pm_word14,pm_word13,pm_word12,pm_word11,pm_word10,pm_word9,pm_word8,pm_word7,pm_word6,pm_word5,pm_word4,pm_word3,pm_word2,pm_word1,pm_word0},clk,sel,ld_val_reg,instruction,addbus,databus);
    prgrm_cnt PC(start,clk,mode,databus,sel);

    ALU un(databus,alu_flag,dm_word0,dm_word1,fs_cal,fs_shft,shft_wr,clk,alu_out);

    inst_dec  ID(instruction[15:8],rr,r,rv,pm,ra,rp,nop,beginx);
    
    MOV asmA6(rr[6],clk,ld_val_reg,mode[0],rd,rd_latch,wr);
    AND asmA5(rr[5],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    OR  asmA4(rr[4],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    ADD asmA3(rr[3],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    SUB asmA2(rr[2],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    XOR asmA1(rr[1],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    CMP asmA0(rr[0],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);

    CLR  asmB6(r[6],clk,ld_val_reg,mode[0],clr);
    NEG  asmB5(r[5],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,databus[0],fs_cal,addbus);
    SLL  asmB4(r[4],clk,ld_val_reg,mode[0],rd,rd_latch,wr,shft_wr,alu_write,fs_shft);
    SLR  asmB3(r[3],clk,ld_val_reg,mode[0],rd,rd_latch,wr,shft_wr,alu_write,fs_shft);
    ROL  asmB2(r[2],clk,ld_val_reg,mode[0],rd,rd_latch,wr,shft_wr,alu_write,fs_shft);
    ROR  asmB1(r[1],clk,ld_val_reg,mode[0],rd,rd_latch,wr,shft_wr,alu_write,fs_shft);
    INC  asmB0(r[0],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,databus[0],fs_cal,addbus);

    LDI  asmC4(rv[4],clk,ld_val_reg,mode[0],wr);
    ANDI asmC3(rv[3],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    ORI  asmC2(rv[2],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    ADI  asmC1(rv[1],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    SBI  asmC0(rv[0],clk,ld_val_reg,mode[0],rd,rd_latch,wr,alu_write,fs_cal,addbus);
    
    JMP  asmD3(pm[3],clk,ld_val_reg,mode);
    BREQ asmD2(pm[2],clk,dm_word32[5],ld_val_reg,mode);
    BRZ  asmD1(pm[1],clk,dm_word32[1],ld_val_reg,mode);
    JPRL  asmD0(pm[0],clk,ld_val_reg,mode);

    LDA  asmE1(ra[1],clk,start,ld_val_reg,mode[0],rd,rd_latch,wr,point_add[26],addbus);
    STA  asmE0(ra[0],clk,start,ld_val_reg,mode[0],rd,rd_latch,wr);

    LDP  asmF1(rp[1],clk,instruction[5],ld_val_reg,mode[0],rd,rd_latch,wr,point_add[31:28]);
    STP  asmF0(rp[0],clk,instruction[5],ld_val_reg,mode[0],rd,rd_latch,wr,point_add[31:28]);

    initial begin
        pm_word0=16'b0010000000000000;      //beginx
        pm_word1=16'b0111100000011111;      //clr R31
        pm_word2=16'b1111010001010101;      // ldi r12 $55
        pm_word3=16'b1000101111101100;      //Sub r31 r12       // pm_word4=16'h1000; 
        pm_word4=16'b0100000000001100;      //inc r12
        pm_word5=16'b0111000000001100;      //neg r12
        pm_word6=16'h1000;
        pm_word7=16'b1011101100001100;      //mov r24 r12
        pm_word8=16'b1100110001010110;      //adi r12 $56
        pm_word9=16'b0110000000000000;      //sll r0
       pm_word10=16'h1000;
       pm_word11=16'b1111110010000000;      // jmp 128
      pm_word128=16'h1000;
      pm_word129=16'b1111100010001110;      //jprl 256-129+15
      pm_word15=16'h1000;
      pm_word16=16'b1111011110000000;      //ldi r15 10000000
      pm_word17=16'b1011101111001111;      //mov r30 r15
      pm_word18=16'b1111011100000011;      //ldi r15 00000011
      pm_word19=16'b1011101111101111;      //mov r31 r15
      pm_word20=16'b0111110111101111;      //stp R15 (896-0011100000)
      pm_word21=16'h1000; 
      pm_word22=16'b1011111000010011;      //lda r19 896
      pm_word23=16'b0000001110000000;      //896 
      pm_word24=16'h1000;
    end

    initial begin
        #11 start=1;
        #1 start=0;
        $dumpfile("test.vcd");
        $dumpvars(0,clrtest);
        $monitor($time,"  %b   %b   %b  %b",nop,mode,databus,dm_word32);
        #1000 $finish;
    end
endmodule

